`timescale 1ns / 1ps
`default_nettype none

module image_resize #(parameter WIDTH = 8) (
                    input wire clk_in,
                    input wire rst_in,

                    output logic error_out,
                    output logic busy_out);

endmodule
