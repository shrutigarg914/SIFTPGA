`timescale 1ns / 1ps
`default_nettype none

// receive two images
// pass them through dog
// transmit result to laptop
// NOTE that we can't send 9 bits over tx
// go from 8 bit greyscale to 7 bit greyscale?
// do some voodoo to squeeze resulting image? (add 2**8 and then divide by 2?)
module top_level(
  input wire [15:0] sw, //all 16 input slide switches
  input wire clk_100mhz,
  input wire uart_rxd,
  input wire [3:0] btn, //all four momentary button switches
  output logic [2:0] rgb0, //rgb led
  output logic [2:0] rgb1, //rgb led
  output logic uart_txd,
  output logic [15:0] led //16 green output LEDs (located right above switches)
  );
    //shut up those rgb LEDs (active high):
    assign rgb1= 0;
    assign rgb0 = 0;

    logic sys_rst;
    assign sys_rst = btn[0];

    parameter DIMENSION = 64;

    logic [13:0] pixel_addr;
    logic [7:0] rx_data;

    logic valid_o;
    logic valid_o_edge;
    logic old_valid_o;

    always_ff @(posedge clk_100mhz) begin
      if (valid_o==old_valid_o) begin
        valid_o_edge <= 1'b0;
      end else begin
        old_valid_o <= valid_o;
        valid_o_edge <= valid_o;
      end
    end

    // TODO: receive image sent over via python script
    uart_rx #(.CLOCKS_PER_BAUD(50))
      urx (
        .clk(clk_100mhz),
        .rx(uart_rxd),
        .data_o(rx_data),
        .valid_o(valid_o)
      );
    logic full_image_received;
    assign led[0] = full_image_received;

    // if we have a valid_o, update pixel location for BRAM 
    always_ff @(posedge clk_100mhz) begin
      if (sys_rst) begin
        pixel_addr <= 0;
        full_image_received <= 1'b0;
      end
      else if (valid_o_edge) begin
        pixel_addr <= pixel_addr + 1;
        if (pixel_addr== DIMENSION*DIMENSION - 1) begin
          full_image_received <= 1'b1;
        end
      end else begin
        if (full_image_received & ~old_full_img) begin 
            full_image_received <= 1'b0;
            // switch which BRAM you're writing to
        end
    end
    // the start image BRAM
    xilinx_true_dual_port_read_first_2_clock_ram #(
    .RAM_WIDTH(8), // we expect 8 bit greyscale images
    .RAM_DEPTH(DIMENSION*DIMENSION)) //we expect a 64*64 image with 16384 pixels total
    img_1 (
    .addra(pixel_addr),
    .clka(clk_100mhz),
    .wea(valid_o),
    .dina(rx_data),
    .ena(1'b1),
    .regcea(1'b1),
    .rsta(sys_rst),
    .douta(), //never read from this side
    .addrb(read_pixel_addr),// transformed lookup pixel
    .dinb(),
    .clkb(clk_100mhz),
    .web(1'b0),
    .enb(1'b1),
    .rstb(sys_rst),
    .regceb(1'b1),
    .doutb(pixel_out)
  );
    xilinx_true_dual_port_read_first_2_clock_ram #(
    .RAM_WIDTH(9), // we expect 8 bit greyscale images
    .RAM_DEPTH(DIMENSION*DIMENSION)) //we expect a 64*64 image with 16384 pixels total
    img_1 (
    .addra(pixel_addr),
    .clka(clk_100mhz),
    .wea(valid_o),
    .dina(rx_data),
    .ena(1'b1),
    .regcea(1'b1),
    .rsta(sys_rst),
    .douta(), //never read from this side
    .addrb(read_pixel_addr),// transformed lookup pixel
    .dinb(),
    .clkb(clk_100mhz),
    .web(1'b0),
    .enb(1'b1),
    .rstb(sys_rst),
    .regceb(1'b1),
    .doutb(pixel_out)
  );

    // TODO: when btn[1] pressed, send what's stored in the output BRAM to the laptop
    
    // button press detected by 
    logic btn_edge;

    //rest of the logic here
    logic start_i;
    logic done_o;
    logic [7:0] data_i;
    logic btn_pulse;
    logic old_btn_pulse;
    debouncer btn1_db(.clk_in(clk_100mhz),
                    .rst_in(sys_rst),
                    .dirty_in(btn[1]),
                    .clean_out(btn_pulse));
 
    /* this should go high for one cycle on the
    * rising edge of the (debounced) button output
    */ 
    /* TODO: write your edge detector for part 1 of the
    * lab here!
    */
    always_ff @(posedge clk_100mhz) begin
      if (btn_pulse==old_btn_pulse) begin
        btn_edge <= 1'b0;
      end else begin
        old_btn_pulse <= btn_pulse;
        btn_edge <= btn_pulse;
      end
    end

    send_img  tx_img (
      .clk(clk_100mhz),
      .rst_in(sys_rst),//sys_rst
      .img_ready(btn_edge),//full_image_received
      .tx(uart_txd),//uart_txd
      .data(pixel_out),
      .address(read_pixel_addr), // gets wired to the BRAM
      .tx_free(led[2]),
      // .out_state(led[4:3]),
      .busy(tx_img_busy) //or we could do img_sent whichever makes more sense
    );
  logic tx_img_busy;

  logic [7:0] pixel_out;
  logic [13:0] read_pixel_addr;
  assign led[1] = tx_img_busy;
  assign led[15:3] = read_pixel_addr[12:0];
  
    
endmodule // top_level

`default_nettype wire
